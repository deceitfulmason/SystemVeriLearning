module cnt_127361(



    
)