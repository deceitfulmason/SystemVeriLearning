module top (
    input  logic         CLK50,
    input  logic [17:0]  SW,
    input  logic  [3:0]  KEY,
    output logic [17:0]  LEDR,
    output logic [8:0]   LEDG,
    output logic [6:0]   HEX [7:0]
);
 


 
/*
 maioria maioria0 (
    .A(SW[0]),
    .B(SW[1]),
    .C(SW[2]),
    .X(SW[3]),
    .Y(LEDG[8])


 );
*/



endmodule