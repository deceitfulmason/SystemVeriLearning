module cod16_4 (
    logic input [15:0] X,
    logic output Y,
    logic output GATE
);

    always_comb begin

        


    end



endmodule