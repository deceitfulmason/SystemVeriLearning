module cod16_4 (
    logic input [15:0]  X,
    logic output        Y,
    logic output        GATE
);

    always_comb begin

       Y = 4'b0000 //Initializes Y as a 4 bit value of 0 to avoid errors 

        
    end



endmodule