module d7s(
    input logic [3:0] X ,
    input logic [0] EN ,
    output logic [6:0] Y 



always_comb begin : 
    
        
    

                if (EN)
        begin 


        end

        else begin



        end

end