module div50m(
    input logic CLK_IN,
    output logic CLK_OUT
);


always_ff @(posedge CLK_IN) begin




end



endmodule