module d7s(
    input logic X [3:0],
    input logic EN [0],
    output logic Y [6:0]

        if (EN)
begin 


end

else begin



end