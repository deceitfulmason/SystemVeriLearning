module cntbit(
input logic X,

);





/*
7. Make an 8-bit counter that:
a) Shows the output in hexadecimal on two 7-segment displays, and in binary on
LEDR[7:0].
b) Increments by one when the user presses KEY[0] and releases it in less than
one second.
c) Returns to zero when the user holds KEY[0] for more than one second.
*/